// som_pkg.vh

`ifndef _som_pkg_vh_
`define _som_pkg_vh_

`define PART_NUM_MAJOR  10'd1
`define PART_NUM_MINOR  6'd1

`define FAST_DIV 75
`define SLOW_DIV 75000
`define ONEM_DIV 1000000

`define MAX_TIME 13'd5000
`define MIN_TIME 13'd1000
`define MAX_SUM  17'd5000
`define MIN_SUM  17'd1000
`define MAX_ARC  4'd15
`define MAX_KV   16'h8000

`endif  //_som_pkg_vh_
